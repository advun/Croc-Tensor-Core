package matrix_pkg;

parameter indata_size = 8;

endpackage 